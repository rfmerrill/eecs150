
module MIPS150(
    input clk, rst,
    input FPGA_SERIAL_RX,
    output FPGA_SERIAL_TX
);

// Use this as the top-level module for your CPU. You
// will likely want to break control and datapath out
// into separate modules that you instantiate here.



endmodule
    

