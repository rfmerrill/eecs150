module MemoryStageControl(input [31:0] ALUOut,
                          input [31:0] WriteData,
                          input [4:0] WriteReg,
                          input );

endmodule
