module MemoryUnMap ();
                     

endmodule
