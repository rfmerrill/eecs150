module MemoryStageControl(input clk, input rst);
  always @(*) begin

  end

  always @(posedge clk) begin

  end

endmodule
